pBAV        k       @       �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@            �@             @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               @<          ��               :��h��TD�|z���x�t��X� � 4�����X                                                                                                                                                                                                                                                                                                                                                                                                                                                               